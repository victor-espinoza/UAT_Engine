`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Author:        Victor Espinoza
// Email:         victor.alfonso94@gmail.com
// Project #:     Project 2 - PicoBlaze Integration with Interrupts 
// Course:        CECS 460
// Create Date:   13:19:08 04/18/2015 
//
// Module Name:   top_level
// File Name:     top_level.v 
//
// Description:   This Display Controller module controls the 7-Segment display
//                and everything that it needs in order to correctly display
//                the appropriate values. This module was created in Professor
//                Allison's CECS 301 class. Each section of this module is 
//                described within the module itself using comments.
//
//
// Dependencies:
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module display_controller(clk, rstb, annode3, annode2, annode1, annode0,  
								  a3, a2, a1, a0, a, b, c, d, e, f, g);
   
   //Input and Output Declarations  
   input           clk, rstb;
   input [3:0]     annode3, annode2, annode1, annode0;
   
   //annode and cathode variables for the 7-Segment Display
   output reg     a, b, c, d, e, f, g;
   output wire    a3, a2, a1, a0;
	
   //Local Variables
   reg  [3:0]      ad_out; 
   wire [1:0]      seg_sel;
   reg             clk_250;
   //counter variable
   reg [15:0]      count = 0;
	
   //initialize LED clock:
   //Divide 50MHz on-board clock to 250Hz. This is done so that
   //it appears to the human observer that all four anode signals
   //are on even when in reality they are not. This is done by
   //driving the cathode patterns at least once every 16ms,
   //which comes out to 4ms per annode/cathode pattern.			  
   always @(posedge clk, negedge rstb)
      //if rstb then rstb count and clock
      if(!rstb) begin
         count <= 0;
         clk_250 <= 0;
      end 
      else begin
         //increment count
         count <= (count + 1);
         //set output clock to opposite if count is greater than or equal to 25000
         if(count >= 25000) begin
            count <= 0;
            clk_250 <= ~clk_250;
         end 
      end
	
	
   //initialize LED controller module:
   //module led_controller(clk, rstb, a3, a2, a1, a0, seg_sel);
   led_controller LED_contr(
	   .clk(clk_250), 
      .rstb(rstb), 
      .a3(a3), 
      .a2(a2), 
      .a1(a1), 
      .a0(a0), 
      .seg_sel(seg_sel)
   );
   
	
   //initialize address mux:
   //This multiplexer is used to select what data input is to 
   //be assigned to the ad_out output and driven to the seven segment
   //display. The value of the ad_out is chosen based on the seg_sel
   //input that was generated by our led_controller module.
   always @(seg_sel, annode3, annode2, annode1, annode0)	
      case (seg_sel)		
         2'b00  :		ad_out =  annode0;  //annode 0
         2'b01  :		ad_out =  annode1;  //annode 1
         2'b10  :		ad_out =  annode2;  //annode 2
         2'b11  :		ad_out =  annode3;  //annode 3
         default: 	ad_out =  4'bx;  //default output	
      endcase		
	

   //initialize hex to seven segment display 
   //This hex_to_7segment module basicaly takes in a four bit input
   //and depending on what that input is, it then transfers that 
   //information by turning on the appropriate segments (a-g) on the 
   //seven segment display in order to represent that four bit input.
   //This was achieved by using case statements for all of the 
   //appropriate 4-bit input options and assigning the according
   //values for a-g for that 4-bit input. Depending on the 4-bit
   //value, the appropriate segments are turned on in order to 
   //display that value.
   always@(ad_out)
      case (ad_out)
         4'b0000: {a, b, c, d, e, f, g} = 7'b0000001; //Display 0
         4'b0001: {a, b, c, d, e, f, g} = 7'b1001111; //Display 1
         4'b0010: {a, b, c, d, e, f, g} = 7'b0010010; //Display 2
         4'b0011: {a, b, c, d, e, f, g} = 7'b0000110; //Display 3
         4'b0100: {a, b, c, d, e, f, g} = 7'b1001100; //Display 4
         4'b0101: {a, b, c, d, e, f, g} = 7'b0100100; //Display 5
         4'b0110: {a, b, c, d, e, f, g} = 7'b0100000; //Display 6
         4'b0111: {a, b, c, d, e, f, g} = 7'b0001111; //Display 7
         4'b1000: {a, b, c, d, e, f, g} = 7'b0000000; //Display 8
         4'b1001: {a, b, c, d, e, f, g} = 7'b0001100; //Display 9
         4'b1010: {a, b, c, d, e, f, g} = 7'b0001000; //Display A
         4'b1011: {a, b, c, d, e, f, g} = 7'b1100000; //Display B
         4'b1100: {a, b, c, d, e, f, g} = 7'b0110001; //Display C
         4'b1101: {a, b, c, d, e, f, g} = 7'b1000010; //Display D
         4'b1110: {a, b, c, d, e, f, g} = 7'b0110000; //Display E
         4'b1111: {a, b, c, d, e, f, g} = 7'b0111000; //Display F
         default: {a, b, c, d, e, f, g} = 7'b1111111; //Display Nothing
      endcase

endmodule
